library ieee;
use ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;

entity instrMemory is
  port (
    Addr: in std_logic_vector(3 downto 0);
    Instruction: out std_logic_vector(31 downto 0)
  );
end instrMemory;

architecture arch1 of instrMemory is

type instr_array is array (0 to 15) of std_logic_vector (31 downto 0);
constant instrmem: instr_array := (
  "00000000010001100010000000100000", -- add $4,$2,$6
  "00000000010001100010100000100010", -- sub $5,$2,$6
  "00000000101001000011000000100000", -- add $6,$5,$4
  "00000000000000000000000000000000",
  "11111111111111111111111111111111",
  "11111111111111111111111111111111",
  "00000000101001100010000000100000", -- add $4,$5,$6
  "11111111111111111111111111111111",
  "11111111111111111111111111111111",
  "11111111111111111111111111111111",
  "11111111111111111111111111111111",
  "11111111111111111111111111111111",
  "11111111111111111111111111111111",
  "11111111111111111111111111111111",
  "11111111111111111111111111111111",
  "11111111111111111111111111111111"
);

begin

  Instruction <= instrmem(to_integer(unsigned(Addr)));

end arch1;
